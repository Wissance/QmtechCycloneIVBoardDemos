

module serial_echo();
endmodule
